/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2021-04-03 13:35:39 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module tb_test_top_sim();
//==========================================================================
//-------- define ----------------------------------------------------------
string test_unit_region;
logic [0-1:0]  unit_pass_u ;
logic [0-1:0]  unit_pass_d ;

//==========================================================================
//-------- instance --------------------------------------------------------
test_top_sim rtl_top(
/* input clock */.sys_clock ( ),
/* output      */.odata     ( )
);
//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
