/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2021-04-03 12:04:33 +0800
madified:
***********************************************/


package head_package;
parameter  HDSIZE = 8;
//==========================================================================
//-------- define ----------------------------------------------------------
typedef struct {
logic [4-1:0]  idata ;
logic valid;
} s_head;


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endpackage:head_package
