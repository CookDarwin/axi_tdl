/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2021-03-20 12:10:27 +0800
madified:
***********************************************/


module test_packageparameter  NUM = 6;();
//==========================================================================
//-------- define ----------------------------------------------------------
typedef struct {
logic [32-1:0]  op ;
logic [NUM-1:0]  pl ;
} s_ing;

typedef struct {
logic [32-1:0]  op ;
logic [NUM-1:0]  pl ;
} z_ing;

logic [32-1:0]  data ;
z_ing zing_v0;
s_ing s_ing_v1;

//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------
assign zing_v0.op[9] = 0;

endmodule
