package SystemPkg;
    parameter SIM = "ON";

endpackage