/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2023-02-17 21:27:53 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module test_top (
    input             sys_clock,
    output logic[3:0] odata
);

//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
