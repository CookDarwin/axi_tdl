/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2021-04-03 13:14:02 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module example_pkg import head_package::*;(
    input [HDSIZE-1:0] indata,
    output logic[31:0] odata
);

//------>> EX CODE <<-------------------
import body_package::*;
//------<< EX CODE >>-------------------

//==========================================================================
//-------- define ----------------------------------------------------------
logic [BDSIZE-1:0]  gdata ;
s_head ss_head;

//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------
assign ss_head.idata = 4;
assign ss_head.valid = 1'b1;

endmodule
