/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2021-03-20 12:10:27 +0800
madified:
***********************************************/


module head_packageparameter  HDSIZE = 8;();
//==========================================================================
//-------- define ----------------------------------------------------------
typedef struct {
logic [4-1:0]  idata ;
logic valid;
} s_head;


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
