/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2025-12-12 04:47:03 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module test_top (
    input             sys_clock,
    output logic[3:0] odata
);

//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
