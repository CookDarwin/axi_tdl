/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2021-03-20 12:10:27 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module tb_test_top();
//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------
test_top rtl_top(
/* input clock */.sys_clock ( ),
/* output      */.odata     ( )
);
//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
