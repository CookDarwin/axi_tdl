package SystemPkg;
    parameter SIM = "OFF";

endpackage