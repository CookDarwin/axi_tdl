/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2022-07-10 11:18:28 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module tb_exp_test_unit_sim();
//==========================================================================
//-------- define ----------------------------------------------------------
logic  sys_clk;
string test_unit_region;
logic [0-1:0]  unit_pass_u ;
logic [0-1:0]  unit_pass_d ;

//==========================================================================
//-------- instance --------------------------------------------------------
exp_test_unit_sim rtl_top(
/* input clock */.clock (sys_clk ),
/* input reset */.rst_n (1'b1    )
);
//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
