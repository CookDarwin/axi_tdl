/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2023-02-17 21:27:54 +0800
madified:
***********************************************/
`timescale 1ns/1ps
`include "define_macro.sv" 

module test_vcs_string #(
    `parameter_longstring(111) INIT_FILE = "ppppppppp"
)();
//==========================================================================
//-------- define ----------------------------------------------------------


//==========================================================================
//-------- instance --------------------------------------------------------

//==========================================================================
//-------- expression ------------------------------------------------------

endmodule
