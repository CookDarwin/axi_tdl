/**********************************************
_______________________________________ 
___________    Cook Darwin   __________    
_______________________________________
descript:
author : Cook.Darwin
Version: VERA.0.0
created: 2021-03-20 20:34:51 +0800
madified:
***********************************************/
`timescale 1ns/1ps

module tb_test_top();
//==========================================================================
//-------- define ----------------------------------------------------------
logic gl_clk;

//==========================================================================
//-------- instance --------------------------------------------------------
test_top rtl_top(
/* input clock */.global_sys_clk (gl_clk )
);
//==========================================================================
//-------- expression ------------------------------------------------------
initial begin
    forever begin #(33ns);gl_clk = ~gl_clk;end;
end

endmodule
